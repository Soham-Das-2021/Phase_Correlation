//*** Design to convert decimal nos.(Image data) into 32 bit Single Precision Floating Point binary nos.
//Conversion happens through the test bench

module test_design_16x16 (clk );
input clk;
reg b;
reg a;

always@(posedge clk)
a =b;

endmodule
